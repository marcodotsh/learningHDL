package barrelshifter_pkg;
  parameter int W = 5;
endpackage
