package barrelshifter_pkg;
  parameter int W = 6;
endpackage
