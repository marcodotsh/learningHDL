package flipflop_pkg;
  parameter int W = 2;
endpackage
