package rrprioassign_pkg;
  parameter int N = 8;
endpackage
